`timescale 1ns/1ns
module mux2_to_1 (input a,b,s,en,output w);
	wire i,j;
	notif1 #(14,18,16) n1(i,a,j);
	notif1 #(14,18,16) n2(i,b,s);
	not #(7,9) n3(j,s);
	notif1 #(14,18,16) n4(w,i,en);
endmodule
module D_latch(input d,clk,en,output q);
	mux2_to_1 mx(q,d,clk,en,q);
endmodule
module ms_DFF(input d,clk,reset,en,output q);
	wire i,j,k,d2,q1;
	not #(7,9) n1(i,reset);
	not #(7,9) n2(j,clk);
	nand #(14,10) o1(k,i,q1);
	not #(7,9) n3(d2,k);
	D_latch dl1(d,clk,en,q1);
	D_latch dl2(d2,j,en,q);
endmodule
module register8withMSDFF(input serIn,clk,reset,en,output [7:0] po);
	wire [8:0] d;
	assign d[8]=serIn;
	genvar k;
	generate
		for(k=8;k>0;k=k-1) begin : registerGates
			ms_DFF dd(d[k],clk,reset,en,d[k-1]);
		end
	endgenerate
	assign po=d[7:0];
endmodule
module register8withAlways(input serIn,clk,reset,en,output logic [7:0] po);
	always @(posedge clk) begin
		if(reset)
			#50 po<=8'b0;
		else 
			#50 po<={serIn,po[7:1]};
	end
endmodule

