`timescale 1ns/1ns
module ALU1 (input signed [15:0] inM,inN,input [2:0] opc,input inC,output zer,neg,output logic signed [15:0] outF);
	assign zer=~(|outF);
	assign neg=outF[15];
	always @(inM,inN,opc,inC) begin
		outF=16'd0;
		case(opc)
			3'd0:outF=inM+inN+inC;
			3'd1:outF=inM+(inN>>>1);
			3'd2:outF=inM+1;
			3'd3:outF=inM+(inM>>>1);
			3'd4:outF=inM&inN;
			3'd5:outF=inM|inN;
			3'd6:outF=~inM;
			3'd7:outF=16'd0;
			default:outF=16'd0;
		endcase
	end
endmodule


module NOT(A, Y);
input A;
output Y;
assign Y = ~A;
endmodule

module NAND(A, B, Y);
input A, B;
output Y;
assign Y = ~(A & B);
endmodule

module NOR(A, B, Y);
input A, B;
output Y;
assign Y = ~(A | B);
endmodule

module DFF(C, D, Q);
input C, D;
output logic Q;
always @(posedge C)
	Q <= D;
endmodule



module ALU2(inM, inN, opc, inC, zer, neg, outF);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  input inC;
  input [15:0] inM;
  input [15:0] inN;
  output neg;
  input [2:0] opc;
  output [15:0] outF;
  output zer;
  NOR _1310_ (
    .A(_0460_),
    .B(_0459_),
    .Y(_0934_)
  );
  NOT _1311_ (
    .A(_0459_),
    .Y(_0945_)
  );
  NOT _1312_ (
    .A(_0460_),
    .Y(_0956_)
  );
  NOR _1313_ (
    .A(_0956_),
    .B(_0945_),
    .Y(_0966_)
  );
  NOR _1314_ (
    .A(_0966_),
    .B(_0934_),
    .Y(_0977_)
  );
  NOT _1315_ (
    .A(_0674_),
    .Y(_0988_)
  );
  NOT _1316_ (
    .A(_0783_),
    .Y(_0998_)
  );
  NOR _1317_ (
    .A(_0998_),
    .B(_0988_),
    .Y(_1019_)
  );
  NOT _1318_ (
    .A(_1019_),
    .Y(_1031_)
  );
  NOR _1319_ (
    .A(_0783_),
    .B(_0674_),
    .Y(_1032_)
  );
  NOR _1320_ (
    .A(_1032_),
    .B(_1019_),
    .Y(_1053_)
  );
  NOT _1321_ (
    .A(_1295_),
    .Y(_1065_)
  );
  NOT _1322_ (
    .A(_1297_),
    .Y(_1066_)
  );
  NOR _1323_ (
    .A(_1066_),
    .B(_1065_),
    .Y(_1077_)
  );
  NOT _1324_ (
    .A(_1077_),
    .Y(_1098_)
  );
  NOR _1325_ (
    .A(_1297_),
    .B(_1295_),
    .Y(_1110_)
  );
  NOT _1326_ (
    .A(_1110_),
    .Y(_1112_)
  );
  NOT _1327_ (
    .A(_1300_),
    .Y(_1133_)
  );
  NOT _1328_ (
    .A(_1302_),
    .Y(_1145_)
  );
  NOR _1329_ (
    .A(_1145_),
    .B(_1133_),
    .Y(_1146_)
  );
  NOT _1330_ (
    .A(_1146_),
    .Y(_1156_)
  );
  NOR _1331_ (
    .A(_1302_),
    .B(_1300_),
    .Y(_1167_)
  );
  NOR _1332_ (
    .A(_1167_),
    .B(_1146_),
    .Y(_1177_)
  );
  NOT _1333_ (
    .A(_1009_),
    .Y(_1188_)
  );
  NOT _1334_ (
    .A(_1020_),
    .Y(_1199_)
  );
  NOR _1335_ (
    .A(_1199_),
    .B(_1188_),
    .Y(_1209_)
  );
  NOT _1336_ (
    .A(_1209_),
    .Y(_1221_)
  );
  NOR _1337_ (
    .A(_1020_),
    .B(_1009_),
    .Y(_1232_)
  );
  NOT _1338_ (
    .A(_1232_),
    .Y(_1242_)
  );
  NOT _1339_ (
    .A(_1043_),
    .Y(_1253_)
  );
  NOT _1340_ (
    .A(_1054_),
    .Y(_1263_)
  );
  NOR _1341_ (
    .A(_1263_),
    .B(_1253_),
    .Y(_1273_)
  );
  NOT _1342_ (
    .A(_1273_),
    .Y(_1284_)
  );
  NOR _1343_ (
    .A(_1054_),
    .B(_1043_),
    .Y(_1293_)
  );
  NOR _1344_ (
    .A(_1293_),
    .B(_1273_),
    .Y(_1294_)
  );
  NOR _1345_ (
    .A(_1099_),
    .B(_1087_),
    .Y(_1296_)
  );
  NOT _1346_ (
    .A(_1087_),
    .Y(_1298_)
  );
  NOT _1347_ (
    .A(_1099_),
    .Y(_1299_)
  );
  NOR _1348_ (
    .A(_1299_),
    .B(_1298_),
    .Y(_1301_)
  );
  NOT _1349_ (
    .A(_1122_),
    .Y(_1303_)
  );
  NOT _1350_ (
    .A(_1134_),
    .Y(_1304_)
  );
  NOR _1351_ (
    .A(_1304_),
    .B(_1303_),
    .Y(_1305_)
  );
  NOT _1352_ (
    .A(_1305_),
    .Y(_1306_)
  );
  NOR _1353_ (
    .A(_1134_),
    .B(_1122_),
    .Y(_1307_)
  );
  NOR _1354_ (
    .A(_1307_),
    .B(_1305_),
    .Y(_1308_)
  );
  NOR _1355_ (
    .A(_0729_),
    .B(_0717_),
    .Y(_1309_)
  );
  NOT _1356_ (
    .A(_0717_),
    .Y(_0461_)
  );
  NOT _1357_ (
    .A(_0729_),
    .Y(_0462_)
  );
  NOR _1358_ (
    .A(_0462_),
    .B(_0461_),
    .Y(_0463_)
  );
  NOT _1359_ (
    .A(_0751_),
    .Y(_0464_)
  );
  NOT _1360_ (
    .A(_0762_),
    .Y(_0465_)
  );
  NOR _1361_ (
    .A(_0465_),
    .B(_0464_),
    .Y(_0467_)
  );
  NOT _1362_ (
    .A(_0467_),
    .Y(_0468_)
  );
  NOR _1363_ (
    .A(_0762_),
    .B(_0751_),
    .Y(_0470_)
  );
  NOR _1364_ (
    .A(_0470_),
    .B(_0467_),
    .Y(_0472_)
  );
  NOR _1365_ (
    .A(_0807_),
    .B(_0795_),
    .Y(_0473_)
  );
  NOT _1366_ (
    .A(_0795_),
    .Y(_0475_)
  );
  NOT _1367_ (
    .A(_0807_),
    .Y(_0476_)
  );
  NOR _1368_ (
    .A(_0476_),
    .B(_0475_),
    .Y(_0477_)
  );
  NOT _1369_ (
    .A(_0829_),
    .Y(_0478_)
  );
  NOT _1370_ (
    .A(_0841_),
    .Y(_0479_)
  );
  NOR _1371_ (
    .A(_0479_),
    .B(_0478_),
    .Y(_0480_)
  );
  NOT _1372_ (
    .A(_0480_),
    .Y(_0481_)
  );
  NOR _1373_ (
    .A(_0841_),
    .B(_0829_),
    .Y(_0482_)
  );
  NOR _1374_ (
    .A(_0482_),
    .B(_0480_),
    .Y(_0483_)
  );
  NOT _1375_ (
    .A(_0557_),
    .Y(_0484_)
  );
  NOT _1376_ (
    .A(_0568_),
    .Y(_0486_)
  );
  NOR _1377_ (
    .A(_0486_),
    .B(_0484_),
    .Y(_0487_)
  );
  NOT _1378_ (
    .A(_0487_),
    .Y(_0488_)
  );
  NOR _1379_ (
    .A(_0568_),
    .B(_0557_),
    .Y(_0489_)
  );
  NOT _1380_ (
    .A(_0489_),
    .Y(_0490_)
  );
  NOT _1381_ (
    .A(_0589_),
    .Y(_0491_)
  );
  NOT _1382_ (
    .A(_0600_),
    .Y(_0492_)
  );
  NOR _1383_ (
    .A(_0492_),
    .B(_0491_),
    .Y(_0493_)
  );
  NOT _1384_ (
    .A(_0493_),
    .Y(_0494_)
  );
  NOR _1385_ (
    .A(_0600_),
    .B(_0589_),
    .Y(_0495_)
  );
  NOR _1386_ (
    .A(_0495_),
    .B(_0493_),
    .Y(_0496_)
  );
  NOT _1387_ (
    .A(_1111_),
    .Y(_0497_)
  );
  NOT _1388_ (
    .A(_1220_),
    .Y(_0498_)
  );
  NOR _1389_ (
    .A(_0498_),
    .B(_0497_),
    .Y(_0499_)
  );
  NOT _1390_ (
    .A(_0499_),
    .Y(_0500_)
  );
  NAND _1391_ (
    .A(_0485_),
    .B(_0474_),
    .Y(_0501_)
  );
  NOT _1392_ (
    .A(_0474_),
    .Y(_0502_)
  );
  NOT _1393_ (
    .A(_0485_),
    .Y(_0503_)
  );
  NOR _1394_ (
    .A(_0503_),
    .B(_0502_),
    .Y(_0504_)
  );
  NOR _1395_ (
    .A(_0485_),
    .B(_0474_),
    .Y(_0505_)
  );
  NOR _1396_ (
    .A(_0505_),
    .B(_0504_),
    .Y(_0506_)
  );
  NAND _1397_ (
    .A(_0506_),
    .B(_0516_),
    .Y(_0507_)
  );
  NAND _1398_ (
    .A(_0507_),
    .B(_0501_),
    .Y(_0508_)
  );
  NOR _1399_ (
    .A(_1220_),
    .B(_1111_),
    .Y(_0509_)
  );
  NOR _1400_ (
    .A(_0509_),
    .B(_0499_),
    .Y(_0510_)
  );
  NAND _1401_ (
    .A(_0510_),
    .B(_0508_),
    .Y(_0511_)
  );
  NAND _1402_ (
    .A(_0511_),
    .B(_0500_),
    .Y(_0512_)
  );
  NAND _1403_ (
    .A(_0512_),
    .B(_0496_),
    .Y(_0513_)
  );
  NAND _1404_ (
    .A(_0513_),
    .B(_0494_),
    .Y(_0514_)
  );
  NAND _1405_ (
    .A(_0514_),
    .B(_0490_),
    .Y(_0515_)
  );
  NAND _1406_ (
    .A(_0515_),
    .B(_0488_),
    .Y(_0517_)
  );
  NAND _1407_ (
    .A(_0517_),
    .B(_0483_),
    .Y(_0518_)
  );
  NAND _1408_ (
    .A(_0518_),
    .B(_0481_),
    .Y(_0519_)
  );
  NOR _1409_ (
    .A(_0519_),
    .B(_0477_),
    .Y(_0520_)
  );
  NOR _1410_ (
    .A(_0520_),
    .B(_0473_),
    .Y(_0521_)
  );
  NAND _1411_ (
    .A(_0521_),
    .B(_0472_),
    .Y(_0522_)
  );
  NAND _1412_ (
    .A(_0522_),
    .B(_0468_),
    .Y(_0523_)
  );
  NOR _1413_ (
    .A(_0523_),
    .B(_0463_),
    .Y(_0524_)
  );
  NOR _1414_ (
    .A(_0524_),
    .B(_1309_),
    .Y(_0525_)
  );
  NAND _1415_ (
    .A(_0525_),
    .B(_1308_),
    .Y(_0526_)
  );
  NAND _1416_ (
    .A(_0526_),
    .B(_1306_),
    .Y(_0527_)
  );
  NOR _1417_ (
    .A(_0527_),
    .B(_1301_),
    .Y(_0528_)
  );
  NOR _1418_ (
    .A(_0528_),
    .B(_1296_),
    .Y(_0529_)
  );
  NAND _1419_ (
    .A(_0529_),
    .B(_1294_),
    .Y(_0530_)
  );
  NAND _1420_ (
    .A(_0530_),
    .B(_1284_),
    .Y(_0531_)
  );
  NAND _1421_ (
    .A(_0531_),
    .B(_1242_),
    .Y(_0532_)
  );
  NAND _1422_ (
    .A(_0532_),
    .B(_1221_),
    .Y(_0533_)
  );
  NAND _1423_ (
    .A(_0533_),
    .B(_1177_),
    .Y(_0534_)
  );
  NAND _1424_ (
    .A(_0534_),
    .B(_1156_),
    .Y(_0535_)
  );
  NAND _1425_ (
    .A(_0535_),
    .B(_1112_),
    .Y(_0536_)
  );
  NAND _1426_ (
    .A(_0536_),
    .B(_1098_),
    .Y(_0537_)
  );
  NAND _1427_ (
    .A(_0537_),
    .B(_1053_),
    .Y(_0538_)
  );
  NAND _1428_ (
    .A(_0538_),
    .B(_1031_),
    .Y(_0539_)
  );
  NAND _1429_ (
    .A(_0539_),
    .B(_0977_),
    .Y(_0540_)
  );
  NOR _1430_ (
    .A(_0471_),
    .B(_0469_),
    .Y(_0541_)
  );
  NOT _1431_ (
    .A(_0541_),
    .Y(_0542_)
  );
  NOR _1432_ (
    .A(_0542_),
    .B(_0466_),
    .Y(_0543_)
  );
  NOT _1433_ (
    .A(_0543_),
    .Y(_0544_)
  );
  NOR _1434_ (
    .A(_0539_),
    .B(_0977_),
    .Y(_0545_)
  );
  NOR _1435_ (
    .A(_0545_),
    .B(_0544_),
    .Y(_0546_)
  );
  NAND _1436_ (
    .A(_0546_),
    .B(_0540_),
    .Y(_0547_)
  );
  NOR _1437_ (
    .A(_0998_),
    .B(_0945_),
    .Y(_0548_)
  );
  NOT _1438_ (
    .A(_0548_),
    .Y(_0549_)
  );
  NOR _1439_ (
    .A(_0783_),
    .B(_0459_),
    .Y(_0550_)
  );
  NOR _1440_ (
    .A(_0550_),
    .B(_0548_),
    .Y(_0551_)
  );
  NOR _1441_ (
    .A(_1066_),
    .B(_0988_),
    .Y(_0552_)
  );
  NOT _1442_ (
    .A(_0552_),
    .Y(_0553_)
  );
  NOR _1443_ (
    .A(_1297_),
    .B(_0674_),
    .Y(_0554_)
  );
  NOT _1444_ (
    .A(_0554_),
    .Y(_0555_)
  );
  NOR _1445_ (
    .A(_1145_),
    .B(_1065_),
    .Y(_0556_)
  );
  NOT _1446_ (
    .A(_0556_),
    .Y(_0558_)
  );
  NOR _1447_ (
    .A(_1302_),
    .B(_1295_),
    .Y(_0559_)
  );
  NOR _1448_ (
    .A(_0559_),
    .B(_0556_),
    .Y(_0560_)
  );
  NOR _1449_ (
    .A(_1133_),
    .B(_1199_),
    .Y(_0561_)
  );
  NOT _1450_ (
    .A(_0561_),
    .Y(_0562_)
  );
  NOR _1451_ (
    .A(_1300_),
    .B(_1020_),
    .Y(_0563_)
  );
  NOT _1452_ (
    .A(_0563_),
    .Y(_0564_)
  );
  NOR _1453_ (
    .A(_1263_),
    .B(_1188_),
    .Y(_0565_)
  );
  NOT _1454_ (
    .A(_0565_),
    .Y(_0566_)
  );
  NOR _1455_ (
    .A(_1054_),
    .B(_1009_),
    .Y(_0567_)
  );
  NOR _1456_ (
    .A(_0567_),
    .B(_0565_),
    .Y(_0569_)
  );
  NOR _1457_ (
    .A(_1299_),
    .B(_1253_),
    .Y(_0570_)
  );
  NOT _1458_ (
    .A(_0570_),
    .Y(_0571_)
  );
  NOR _1459_ (
    .A(_1099_),
    .B(_1043_),
    .Y(_0572_)
  );
  NOT _1460_ (
    .A(_0572_),
    .Y(_0573_)
  );
  NOR _1461_ (
    .A(_1304_),
    .B(_1298_),
    .Y(_0574_)
  );
  NOT _1462_ (
    .A(_0574_),
    .Y(_0575_)
  );
  NOR _1463_ (
    .A(_1134_),
    .B(_1087_),
    .Y(_0576_)
  );
  NOR _1464_ (
    .A(_0576_),
    .B(_0574_),
    .Y(_0577_)
  );
  NOR _1465_ (
    .A(_1303_),
    .B(_0462_),
    .Y(_0578_)
  );
  NOT _1466_ (
    .A(_0578_),
    .Y(_0579_)
  );
  NOR _1467_ (
    .A(_1122_),
    .B(_0729_),
    .Y(_0580_)
  );
  NOT _1468_ (
    .A(_0580_),
    .Y(_0581_)
  );
  NOR _1469_ (
    .A(_0465_),
    .B(_0461_),
    .Y(_0582_)
  );
  NOT _1470_ (
    .A(_0582_),
    .Y(_0583_)
  );
  NOR _1471_ (
    .A(_0762_),
    .B(_0717_),
    .Y(_0584_)
  );
  NOR _1472_ (
    .A(_0584_),
    .B(_0582_),
    .Y(_0585_)
  );
  NOR _1473_ (
    .A(_0476_),
    .B(_0464_),
    .Y(_0586_)
  );
  NOT _1474_ (
    .A(_0586_),
    .Y(_0587_)
  );
  NOR _1475_ (
    .A(_0807_),
    .B(_0751_),
    .Y(_0588_)
  );
  NOT _1476_ (
    .A(_0588_),
    .Y(_0590_)
  );
  NOR _1477_ (
    .A(_0479_),
    .B(_0475_),
    .Y(_0591_)
  );
  NOT _1478_ (
    .A(_0591_),
    .Y(_0592_)
  );
  NOR _1479_ (
    .A(_0841_),
    .B(_0795_),
    .Y(_0593_)
  );
  NOR _1480_ (
    .A(_0593_),
    .B(_0591_),
    .Y(_0594_)
  );
  NOR _1481_ (
    .A(_0478_),
    .B(_0486_),
    .Y(_0595_)
  );
  NOT _1482_ (
    .A(_0595_),
    .Y(_0596_)
  );
  NOR _1483_ (
    .A(_0492_),
    .B(_0484_),
    .Y(_0597_)
  );
  NOT _1484_ (
    .A(_0597_),
    .Y(_0598_)
  );
  NOR _1485_ (
    .A(_0491_),
    .B(_0498_),
    .Y(_0599_)
  );
  NOT _1486_ (
    .A(_0599_),
    .Y(_0601_)
  );
  NOR _1487_ (
    .A(_0503_),
    .B(_0497_),
    .Y(_0602_)
  );
  NOR _1488_ (
    .A(_0589_),
    .B(_1220_),
    .Y(_0603_)
  );
  NOR _1489_ (
    .A(_0603_),
    .B(_0599_),
    .Y(_0604_)
  );
  NAND _1490_ (
    .A(_0604_),
    .B(_0602_),
    .Y(_0605_)
  );
  NAND _1491_ (
    .A(_0605_),
    .B(_0601_),
    .Y(_0606_)
  );
  NOR _1492_ (
    .A(_0600_),
    .B(_0557_),
    .Y(_0607_)
  );
  NOR _1493_ (
    .A(_0607_),
    .B(_0597_),
    .Y(_0608_)
  );
  NAND _1494_ (
    .A(_0608_),
    .B(_0606_),
    .Y(_0609_)
  );
  NAND _1495_ (
    .A(_0609_),
    .B(_0598_),
    .Y(_0610_)
  );
  NOR _1496_ (
    .A(_0829_),
    .B(_0568_),
    .Y(_0611_)
  );
  NOR _1497_ (
    .A(_0611_),
    .B(_0595_),
    .Y(_0612_)
  );
  NAND _1498_ (
    .A(_0612_),
    .B(_0610_),
    .Y(_0613_)
  );
  NAND _1499_ (
    .A(_0613_),
    .B(_0596_),
    .Y(_0614_)
  );
  NAND _1500_ (
    .A(_0614_),
    .B(_0594_),
    .Y(_0615_)
  );
  NAND _1501_ (
    .A(_0615_),
    .B(_0592_),
    .Y(_0616_)
  );
  NAND _1502_ (
    .A(_0616_),
    .B(_0590_),
    .Y(_0617_)
  );
  NAND _1503_ (
    .A(_0617_),
    .B(_0587_),
    .Y(_0618_)
  );
  NAND _1504_ (
    .A(_0618_),
    .B(_0585_),
    .Y(_0619_)
  );
  NAND _1505_ (
    .A(_0619_),
    .B(_0583_),
    .Y(_0620_)
  );
  NAND _1506_ (
    .A(_0620_),
    .B(_0581_),
    .Y(_0621_)
  );
  NAND _1507_ (
    .A(_0621_),
    .B(_0579_),
    .Y(_0622_)
  );
  NAND _1508_ (
    .A(_0622_),
    .B(_0577_),
    .Y(_0623_)
  );
  NAND _1509_ (
    .A(_0623_),
    .B(_0575_),
    .Y(_0624_)
  );
  NAND _1510_ (
    .A(_0624_),
    .B(_0573_),
    .Y(_0625_)
  );
  NAND _1511_ (
    .A(_0625_),
    .B(_0571_),
    .Y(_0626_)
  );
  NAND _1512_ (
    .A(_0626_),
    .B(_0569_),
    .Y(_0627_)
  );
  NAND _1513_ (
    .A(_0627_),
    .B(_0566_),
    .Y(_0628_)
  );
  NAND _1514_ (
    .A(_0628_),
    .B(_0564_),
    .Y(_0629_)
  );
  NAND _1515_ (
    .A(_0629_),
    .B(_0562_),
    .Y(_0630_)
  );
  NAND _1516_ (
    .A(_0630_),
    .B(_0560_),
    .Y(_0631_)
  );
  NAND _1517_ (
    .A(_0631_),
    .B(_0558_),
    .Y(_0632_)
  );
  NAND _1518_ (
    .A(_0632_),
    .B(_0555_),
    .Y(_0633_)
  );
  NAND _1519_ (
    .A(_0633_),
    .B(_0553_),
    .Y(_0634_)
  );
  NAND _1520_ (
    .A(_0634_),
    .B(_0551_),
    .Y(_0635_)
  );
  NAND _1521_ (
    .A(_0635_),
    .B(_0549_),
    .Y(_0636_)
  );
  NOR _1522_ (
    .A(_0636_),
    .B(_0977_),
    .Y(_0637_)
  );
  NAND _1523_ (
    .A(_0636_),
    .B(_0977_),
    .Y(_0639_)
  );
  NOT _1524_ (
    .A(_0471_),
    .Y(_0640_)
  );
  NOR _1525_ (
    .A(_0640_),
    .B(_0469_),
    .Y(_0641_)
  );
  NOT _1526_ (
    .A(_0641_),
    .Y(_0642_)
  );
  NOR _1527_ (
    .A(_0642_),
    .B(_0466_),
    .Y(_0643_)
  );
  NAND _1528_ (
    .A(_0643_),
    .B(_0639_),
    .Y(_0644_)
  );
  NOR _1529_ (
    .A(_0644_),
    .B(_0637_),
    .Y(_0645_)
  );
  NOR _1530_ (
    .A(_0998_),
    .B(_0956_),
    .Y(_0646_)
  );
  NOT _1531_ (
    .A(_0646_),
    .Y(_0647_)
  );
  NOR _1532_ (
    .A(_0783_),
    .B(_0460_),
    .Y(_0648_)
  );
  NOR _1533_ (
    .A(_0648_),
    .B(_0646_),
    .Y(_0649_)
  );
  NOR _1534_ (
    .A(_1297_),
    .B(_0783_),
    .Y(_0651_)
  );
  NOR _1535_ (
    .A(_1066_),
    .B(_0998_),
    .Y(_0652_)
  );
  NOR _1536_ (
    .A(_1145_),
    .B(_1066_),
    .Y(_0653_)
  );
  NOT _1537_ (
    .A(_0653_),
    .Y(_0654_)
  );
  NOR _1538_ (
    .A(_1302_),
    .B(_1297_),
    .Y(_0655_)
  );
  NOR _1539_ (
    .A(_0655_),
    .B(_0653_),
    .Y(_0656_)
  );
  NOR _1540_ (
    .A(_1263_),
    .B(_1199_),
    .Y(_0657_)
  );
  NOR _1541_ (
    .A(_1054_),
    .B(_1020_),
    .Y(_0658_)
  );
  NOR _1542_ (
    .A(_0658_),
    .B(_0657_),
    .Y(_0659_)
  );
  NOR _1543_ (
    .A(_1145_),
    .B(_1199_),
    .Y(_0660_)
  );
  NOR _1544_ (
    .A(_1302_),
    .B(_1020_),
    .Y(_0661_)
  );
  NOR _1545_ (
    .A(_0661_),
    .B(_0660_),
    .Y(_0662_)
  );
  NAND _1546_ (
    .A(_0662_),
    .B(_0659_),
    .Y(_0663_)
  );
  NOT _1547_ (
    .A(_0663_),
    .Y(_0664_)
  );
  NOR _1548_ (
    .A(_1299_),
    .B(_1263_),
    .Y(_0665_)
  );
  NOR _1549_ (
    .A(_1099_),
    .B(_1054_),
    .Y(_0666_)
  );
  NOR _1550_ (
    .A(_0666_),
    .B(_0665_),
    .Y(_0667_)
  );
  NOT _1551_ (
    .A(_0667_),
    .Y(_0668_)
  );
  NOR _1552_ (
    .A(_1304_),
    .B(_1299_),
    .Y(_0670_)
  );
  NOR _1553_ (
    .A(_1134_),
    .B(_1099_),
    .Y(_0671_)
  );
  NOR _1554_ (
    .A(_0671_),
    .B(_0670_),
    .Y(_0672_)
  );
  NOR _1555_ (
    .A(_0465_),
    .B(_0462_),
    .Y(_0673_)
  );
  NOR _1556_ (
    .A(_0762_),
    .B(_0729_),
    .Y(_0675_)
  );
  NOR _1557_ (
    .A(_0675_),
    .B(_0673_),
    .Y(_0676_)
  );
  NOT _1558_ (
    .A(_0676_),
    .Y(_0677_)
  );
  NOR _1559_ (
    .A(_0476_),
    .B(_0465_),
    .Y(_0678_)
  );
  NOR _1560_ (
    .A(_0807_),
    .B(_0762_),
    .Y(_0679_)
  );
  NOR _1561_ (
    .A(_0479_),
    .B(_0476_),
    .Y(_0680_)
  );
  NOR _1562_ (
    .A(_0841_),
    .B(_0807_),
    .Y(_0681_)
  );
  NOR _1563_ (
    .A(_0681_),
    .B(_0680_),
    .Y(_0682_)
  );
  NOT _1564_ (
    .A(_0682_),
    .Y(_0683_)
  );
  NOR _1565_ (
    .A(_0841_),
    .B(_0568_),
    .Y(_0684_)
  );
  NOR _1566_ (
    .A(_0479_),
    .B(_0486_),
    .Y(_0686_)
  );
  NOR _1567_ (
    .A(_0492_),
    .B(_0486_),
    .Y(_0687_)
  );
  NOR _1568_ (
    .A(_0600_),
    .B(_0568_),
    .Y(_0688_)
  );
  NOR _1569_ (
    .A(_0688_),
    .B(_0687_),
    .Y(_0689_)
  );
  NOT _1570_ (
    .A(_0689_),
    .Y(_0690_)
  );
  NOR _1571_ (
    .A(_0600_),
    .B(_0485_),
    .Y(_0691_)
  );
  NOR _1572_ (
    .A(_0691_),
    .B(_0498_),
    .Y(_0692_)
  );
  NOT _1573_ (
    .A(_0692_),
    .Y(_0693_)
  );
  NOR _1574_ (
    .A(_0693_),
    .B(_0690_),
    .Y(_0694_)
  );
  NOR _1575_ (
    .A(_0694_),
    .B(_0687_),
    .Y(_0695_)
  );
  NOT _1576_ (
    .A(_0695_),
    .Y(_0696_)
  );
  NOR _1577_ (
    .A(_0696_),
    .B(_0686_),
    .Y(_0697_)
  );
  NOR _1578_ (
    .A(_0697_),
    .B(_0684_),
    .Y(_0698_)
  );
  NOT _1579_ (
    .A(_0698_),
    .Y(_0699_)
  );
  NOR _1580_ (
    .A(_0699_),
    .B(_0683_),
    .Y(_0700_)
  );
  NOR _1581_ (
    .A(_0700_),
    .B(_0680_),
    .Y(_0701_)
  );
  NOR _1582_ (
    .A(_0701_),
    .B(_0679_),
    .Y(_0702_)
  );
  NOR _1583_ (
    .A(_0702_),
    .B(_0678_),
    .Y(_0703_)
  );
  NOR _1584_ (
    .A(_0703_),
    .B(_0677_),
    .Y(_0704_)
  );
  NOR _1585_ (
    .A(_1134_),
    .B(_0729_),
    .Y(_0705_)
  );
  NOT _1586_ (
    .A(_0705_),
    .Y(_0706_)
  );
  NAND _1587_ (
    .A(_0706_),
    .B(_0704_),
    .Y(_0707_)
  );
  NOR _1588_ (
    .A(_1304_),
    .B(_0462_),
    .Y(_0708_)
  );
  NOR _1589_ (
    .A(_0708_),
    .B(_0673_),
    .Y(_0709_)
  );
  NAND _1590_ (
    .A(_0709_),
    .B(_0707_),
    .Y(_0710_)
  );
  NAND _1591_ (
    .A(_0710_),
    .B(_0672_),
    .Y(_0711_)
  );
  NOR _1592_ (
    .A(_0711_),
    .B(_0668_),
    .Y(_0713_)
  );
  NAND _1593_ (
    .A(_0713_),
    .B(_0664_),
    .Y(_0714_)
  );
  NOT _1594_ (
    .A(_0660_),
    .Y(_0715_)
  );
  NOR _1595_ (
    .A(_0670_),
    .B(_0665_),
    .Y(_0716_)
  );
  NOR _1596_ (
    .A(_0716_),
    .B(_0663_),
    .Y(_0718_)
  );
  NOR _1597_ (
    .A(_0718_),
    .B(_0657_),
    .Y(_0719_)
  );
  NAND _1598_ (
    .A(_0719_),
    .B(_0715_),
    .Y(_0720_)
  );
  NOT _1599_ (
    .A(_0720_),
    .Y(_0721_)
  );
  NAND _1600_ (
    .A(_0721_),
    .B(_0714_),
    .Y(_0722_)
  );
  NAND _1601_ (
    .A(_0722_),
    .B(_0656_),
    .Y(_0723_)
  );
  NAND _1602_ (
    .A(_0723_),
    .B(_0654_),
    .Y(_0724_)
  );
  NOR _1603_ (
    .A(_0724_),
    .B(_0652_),
    .Y(_0726_)
  );
  NOR _1604_ (
    .A(_0726_),
    .B(_0651_),
    .Y(_0727_)
  );
  NAND _1605_ (
    .A(_0727_),
    .B(_0649_),
    .Y(_0728_)
  );
  NAND _1606_ (
    .A(_0728_),
    .B(_0647_),
    .Y(_0730_)
  );
  NOT _1607_ (
    .A(_0469_),
    .Y(_0731_)
  );
  NOR _1608_ (
    .A(_0731_),
    .B(_0466_),
    .Y(_0732_)
  );
  NAND _1609_ (
    .A(_0732_),
    .B(_0471_),
    .Y(_0733_)
  );
  NOT _1610_ (
    .A(_0733_),
    .Y(_0734_)
  );
  NAND _1611_ (
    .A(_0734_),
    .B(_0730_),
    .Y(_0735_)
  );
  NOT _1612_ (
    .A(_0678_),
    .Y(_0736_)
  );
  NOT _1613_ (
    .A(_0686_),
    .Y(_0737_)
  );
  NOR _1614_ (
    .A(_0503_),
    .B(_0498_),
    .Y(_0738_)
  );
  NOT _1615_ (
    .A(_0738_),
    .Y(_0739_)
  );
  NOR _1616_ (
    .A(_0739_),
    .B(_0492_),
    .Y(_0740_)
  );
  NOT _1617_ (
    .A(_0740_),
    .Y(_0741_)
  );
  NOR _1618_ (
    .A(_0741_),
    .B(_0737_),
    .Y(_0742_)
  );
  NOT _1619_ (
    .A(_0742_),
    .Y(_0743_)
  );
  NOR _1620_ (
    .A(_0743_),
    .B(_0736_),
    .Y(_0744_)
  );
  NAND _1621_ (
    .A(_0744_),
    .B(_0708_),
    .Y(_0746_)
  );
  NOT _1622_ (
    .A(_0746_),
    .Y(_0747_)
  );
  NAND _1623_ (
    .A(_0747_),
    .B(_0665_),
    .Y(_0748_)
  );
  NOR _1624_ (
    .A(_0748_),
    .B(_1199_),
    .Y(_0749_)
  );
  NOT _1625_ (
    .A(_0749_),
    .Y(_0750_)
  );
  NOR _1626_ (
    .A(_0750_),
    .B(_1145_),
    .Y(_0752_)
  );
  NAND _1627_ (
    .A(_0752_),
    .B(_0652_),
    .Y(_0753_)
  );
  NOR _1628_ (
    .A(_0753_),
    .B(_0956_),
    .Y(_0754_)
  );
  NOR _1629_ (
    .A(_0471_),
    .B(_0731_),
    .Y(_0755_)
  );
  NOT _1630_ (
    .A(_0755_),
    .Y(_0756_)
  );
  NOR _1631_ (
    .A(_0756_),
    .B(_0466_),
    .Y(_0757_)
  );
  NAND _1632_ (
    .A(_0753_),
    .B(_0956_),
    .Y(_0758_)
  );
  NAND _1633_ (
    .A(_0758_),
    .B(_0757_),
    .Y(_0759_)
  );
  NOR _1634_ (
    .A(_0759_),
    .B(_0754_),
    .Y(_0760_)
  );
  NOT _1635_ (
    .A(_0466_),
    .Y(_0761_)
  );
  NOR _1636_ (
    .A(_0542_),
    .B(_0761_),
    .Y(_0763_)
  );
  NAND _1637_ (
    .A(_0763_),
    .B(_0966_),
    .Y(_0764_)
  );
  NOR _1638_ (
    .A(_0756_),
    .B(_0761_),
    .Y(_0766_)
  );
  NOT _1639_ (
    .A(_0766_),
    .Y(_0767_)
  );
  NOR _1640_ (
    .A(_0767_),
    .B(_0460_),
    .Y(_0768_)
  );
  NOR _1641_ (
    .A(_0642_),
    .B(_0761_),
    .Y(_0769_)
  );
  NOT _1642_ (
    .A(_0769_),
    .Y(_0770_)
  );
  NOR _1643_ (
    .A(_0770_),
    .B(_0934_),
    .Y(_0771_)
  );
  NOR _1644_ (
    .A(_0771_),
    .B(_0768_),
    .Y(_0772_)
  );
  NAND _1645_ (
    .A(_0772_),
    .B(_0764_),
    .Y(_0773_)
  );
  NOR _1646_ (
    .A(_0773_),
    .B(_0760_),
    .Y(_0774_)
  );
  NAND _1647_ (
    .A(_0774_),
    .B(_0735_),
    .Y(_0775_)
  );
  NOR _1648_ (
    .A(_0775_),
    .B(_0645_),
    .Y(_0776_)
  );
  NAND _1649_ (
    .A(_0776_),
    .B(_0547_),
    .Y(_0638_)
  );
  NOT _1650_ (
    .A(_1053_),
    .Y(_0777_)
  );
  NOT _1651_ (
    .A(_1177_),
    .Y(_0778_)
  );
  NOT _1652_ (
    .A(_1294_),
    .Y(_0779_)
  );
  NOT _1653_ (
    .A(_1308_),
    .Y(_0780_)
  );
  NOT _1654_ (
    .A(_0472_),
    .Y(_0781_)
  );
  NOT _1655_ (
    .A(_0483_),
    .Y(_0782_)
  );
  NOT _1656_ (
    .A(_0496_),
    .Y(_0784_)
  );
  NOT _1657_ (
    .A(_0516_),
    .Y(_0785_)
  );
  NOT _1658_ (
    .A(_0505_),
    .Y(_0786_)
  );
  NAND _1659_ (
    .A(_0786_),
    .B(_0501_),
    .Y(_0787_)
  );
  NOR _1660_ (
    .A(_0787_),
    .B(_0785_),
    .Y(_0788_)
  );
  NOR _1661_ (
    .A(_0788_),
    .B(_0504_),
    .Y(_0789_)
  );
  NOT _1662_ (
    .A(_0510_),
    .Y(_0790_)
  );
  NOR _1663_ (
    .A(_0790_),
    .B(_0789_),
    .Y(_0791_)
  );
  NOR _1664_ (
    .A(_0791_),
    .B(_0499_),
    .Y(_0793_)
  );
  NOR _1665_ (
    .A(_0793_),
    .B(_0784_),
    .Y(_0794_)
  );
  NOR _1666_ (
    .A(_0794_),
    .B(_0493_),
    .Y(_0796_)
  );
  NOR _1667_ (
    .A(_0796_),
    .B(_0489_),
    .Y(_0797_)
  );
  NOR _1668_ (
    .A(_0797_),
    .B(_0487_),
    .Y(_0798_)
  );
  NOR _1669_ (
    .A(_0798_),
    .B(_0782_),
    .Y(_0799_)
  );
  NOR _1670_ (
    .A(_0799_),
    .B(_0480_),
    .Y(_0800_)
  );
  NOR _1671_ (
    .A(_0800_),
    .B(_0473_),
    .Y(_0801_)
  );
  NOR _1672_ (
    .A(_0801_),
    .B(_0477_),
    .Y(_0802_)
  );
  NOR _1673_ (
    .A(_0802_),
    .B(_0781_),
    .Y(_0803_)
  );
  NOR _1674_ (
    .A(_0803_),
    .B(_0467_),
    .Y(_0804_)
  );
  NOR _1675_ (
    .A(_0804_),
    .B(_1309_),
    .Y(_0806_)
  );
  NOR _1676_ (
    .A(_0806_),
    .B(_0463_),
    .Y(_0808_)
  );
  NOR _1677_ (
    .A(_0808_),
    .B(_0780_),
    .Y(_0809_)
  );
  NOR _1678_ (
    .A(_0809_),
    .B(_1305_),
    .Y(_0810_)
  );
  NOR _1679_ (
    .A(_0810_),
    .B(_1296_),
    .Y(_0811_)
  );
  NOR _1680_ (
    .A(_0811_),
    .B(_1301_),
    .Y(_0812_)
  );
  NOR _1681_ (
    .A(_0812_),
    .B(_0779_),
    .Y(_0813_)
  );
  NOR _1682_ (
    .A(_0813_),
    .B(_1273_),
    .Y(_0814_)
  );
  NOR _1683_ (
    .A(_0814_),
    .B(_1232_),
    .Y(_0815_)
  );
  NOR _1684_ (
    .A(_0815_),
    .B(_1209_),
    .Y(_0816_)
  );
  NOR _1685_ (
    .A(_0816_),
    .B(_0778_),
    .Y(_0817_)
  );
  NOR _1686_ (
    .A(_0817_),
    .B(_1146_),
    .Y(_0818_)
  );
  NOR _1687_ (
    .A(_0818_),
    .B(_1110_),
    .Y(_0819_)
  );
  NOR _1688_ (
    .A(_0819_),
    .B(_1077_),
    .Y(_0820_)
  );
  NAND _1689_ (
    .A(_0820_),
    .B(_0777_),
    .Y(_0821_)
  );
  NAND _1690_ (
    .A(_0821_),
    .B(_0538_),
    .Y(_0823_)
  );
  NAND _1691_ (
    .A(_0823_),
    .B(_0543_),
    .Y(_0824_)
  );
  NOT _1692_ (
    .A(_0551_),
    .Y(_0825_)
  );
  NOT _1693_ (
    .A(_0634_),
    .Y(_0826_)
  );
  NAND _1694_ (
    .A(_0826_),
    .B(_0825_),
    .Y(_0827_)
  );
  NOT _1695_ (
    .A(_0635_),
    .Y(_0828_)
  );
  NOT _1696_ (
    .A(_0643_),
    .Y(_0830_)
  );
  NOR _1697_ (
    .A(_0830_),
    .B(_0828_),
    .Y(_0831_)
  );
  NAND _1698_ (
    .A(_0831_),
    .B(_0827_),
    .Y(_0832_)
  );
  NOR _1699_ (
    .A(_0727_),
    .B(_0649_),
    .Y(_0833_)
  );
  NAND _1700_ (
    .A(_0734_),
    .B(_0728_),
    .Y(_0834_)
  );
  NOR _1701_ (
    .A(_0834_),
    .B(_0833_),
    .Y(_0835_)
  );
  NOT _1702_ (
    .A(_0670_),
    .Y(_0837_)
  );
  NAND _1703_ (
    .A(_0744_),
    .B(_0729_),
    .Y(_0838_)
  );
  NOR _1704_ (
    .A(_0838_),
    .B(_0837_),
    .Y(_0839_)
  );
  NOT _1705_ (
    .A(_0839_),
    .Y(_0840_)
  );
  NOR _1706_ (
    .A(_0840_),
    .B(_1263_),
    .Y(_0842_)
  );
  NAND _1707_ (
    .A(_0842_),
    .B(_0660_),
    .Y(_0843_)
  );
  NOR _1708_ (
    .A(_0843_),
    .B(_1066_),
    .Y(_0844_)
  );
  NOR _1709_ (
    .A(_0844_),
    .B(_0783_),
    .Y(_0845_)
  );
  NAND _1710_ (
    .A(_0753_),
    .B(_0757_),
    .Y(_0846_)
  );
  NOR _1711_ (
    .A(_0846_),
    .B(_0845_),
    .Y(_0847_)
  );
  NOT _1712_ (
    .A(_0763_),
    .Y(_0848_)
  );
  NOR _1713_ (
    .A(_0848_),
    .B(_1031_),
    .Y(_0849_)
  );
  NOR _1714_ (
    .A(_0767_),
    .B(_0783_),
    .Y(_0850_)
  );
  NOR _1715_ (
    .A(_0850_),
    .B(_0849_),
    .Y(_0851_)
  );
  NOR _1716_ (
    .A(_0770_),
    .B(_1032_),
    .Y(_0852_)
  );
  NOR _1717_ (
    .A(_0852_),
    .B(_0543_),
    .Y(_0853_)
  );
  NAND _1718_ (
    .A(_0853_),
    .B(_0851_),
    .Y(_0854_)
  );
  NOR _1719_ (
    .A(_0854_),
    .B(_0847_),
    .Y(_0855_)
  );
  NOT _1720_ (
    .A(_0855_),
    .Y(_0857_)
  );
  NOR _1721_ (
    .A(_0857_),
    .B(_0835_),
    .Y(_0858_)
  );
  NAND _1722_ (
    .A(_0858_),
    .B(_0832_),
    .Y(_0859_)
  );
  NAND _1723_ (
    .A(_0859_),
    .B(_0824_),
    .Y(_0860_)
  );
  NOT _1724_ (
    .A(_0860_),
    .Y(_0650_)
  );
  NOR _1725_ (
    .A(_1110_),
    .B(_1077_),
    .Y(_0861_)
  );
  NOT _1726_ (
    .A(_0861_),
    .Y(_0862_)
  );
  NAND _1727_ (
    .A(_0862_),
    .B(_0535_),
    .Y(_0863_)
  );
  NAND _1728_ (
    .A(_0861_),
    .B(_0818_),
    .Y(_0864_)
  );
  NAND _1729_ (
    .A(_0864_),
    .B(_0863_),
    .Y(_0865_)
  );
  NAND _1730_ (
    .A(_0865_),
    .B(_0543_),
    .Y(_0866_)
  );
  NOR _1731_ (
    .A(_0651_),
    .B(_0652_),
    .Y(_0868_)
  );
  NOR _1732_ (
    .A(_0868_),
    .B(_0724_),
    .Y(_0869_)
  );
  NAND _1733_ (
    .A(_0868_),
    .B(_0724_),
    .Y(_0870_)
  );
  NAND _1734_ (
    .A(_0870_),
    .B(_0734_),
    .Y(_0871_)
  );
  NOR _1735_ (
    .A(_0871_),
    .B(_0869_),
    .Y(_0872_)
  );
  NOR _1736_ (
    .A(_0554_),
    .B(_0552_),
    .Y(_0873_)
  );
  NAND _1737_ (
    .A(_0873_),
    .B(_0632_),
    .Y(_0874_)
  );
  NOR _1738_ (
    .A(_0873_),
    .B(_0632_),
    .Y(_0875_)
  );
  NOR _1739_ (
    .A(_0875_),
    .B(_0830_),
    .Y(_0876_)
  );
  NAND _1740_ (
    .A(_0876_),
    .B(_0874_),
    .Y(_0877_)
  );
  NOT _1741_ (
    .A(_0757_),
    .Y(_0878_)
  );
  NOT _1742_ (
    .A(_0844_),
    .Y(_0879_)
  );
  NAND _1743_ (
    .A(_0843_),
    .B(_1066_),
    .Y(_0881_)
  );
  NAND _1744_ (
    .A(_0881_),
    .B(_0879_),
    .Y(_0882_)
  );
  NOR _1745_ (
    .A(_0882_),
    .B(_0878_),
    .Y(_0883_)
  );
  NAND _1746_ (
    .A(_0769_),
    .B(_1112_),
    .Y(_0884_)
  );
  NOR _1747_ (
    .A(_0767_),
    .B(_1297_),
    .Y(_0885_)
  );
  NOR _1748_ (
    .A(_0848_),
    .B(_1098_),
    .Y(_0886_)
  );
  NOR _1749_ (
    .A(_0886_),
    .B(_0885_),
    .Y(_0887_)
  );
  NAND _1750_ (
    .A(_0887_),
    .B(_0884_),
    .Y(_0888_)
  );
  NOR _1751_ (
    .A(_0888_),
    .B(_0883_),
    .Y(_0889_)
  );
  NAND _1752_ (
    .A(_0889_),
    .B(_0877_),
    .Y(_0891_)
  );
  NOR _1753_ (
    .A(_0891_),
    .B(_0872_),
    .Y(_0892_)
  );
  NAND _1754_ (
    .A(_0892_),
    .B(_0866_),
    .Y(_0669_)
  );
  NAND _1755_ (
    .A(_0816_),
    .B(_0778_),
    .Y(_0893_)
  );
  NAND _1756_ (
    .A(_0893_),
    .B(_0534_),
    .Y(_0894_)
  );
  NAND _1757_ (
    .A(_0894_),
    .B(_0543_),
    .Y(_0895_)
  );
  NOR _1758_ (
    .A(_0630_),
    .B(_0560_),
    .Y(_0896_)
  );
  NOT _1759_ (
    .A(_0896_),
    .Y(_0897_)
  );
  NOT _1760_ (
    .A(_0631_),
    .Y(_0898_)
  );
  NOR _1761_ (
    .A(_0830_),
    .B(_0898_),
    .Y(_0899_)
  );
  NAND _1762_ (
    .A(_0899_),
    .B(_0897_),
    .Y(_0900_)
  );
  NOR _1763_ (
    .A(_0722_),
    .B(_0656_),
    .Y(_0901_)
  );
  NAND _1764_ (
    .A(_0734_),
    .B(_0723_),
    .Y(_0902_)
  );
  NOR _1765_ (
    .A(_0902_),
    .B(_0901_),
    .Y(_0903_)
  );
  NOT _1766_ (
    .A(_0843_),
    .Y(_0904_)
  );
  NOR _1767_ (
    .A(_0749_),
    .B(_1302_),
    .Y(_0906_)
  );
  NOT _1768_ (
    .A(_0906_),
    .Y(_0907_)
  );
  NAND _1769_ (
    .A(_0907_),
    .B(_0757_),
    .Y(_0908_)
  );
  NOR _1770_ (
    .A(_0908_),
    .B(_0904_),
    .Y(_0909_)
  );
  NOR _1771_ (
    .A(_0542_),
    .B(_1156_),
    .Y(_0910_)
  );
  NOR _1772_ (
    .A(_0770_),
    .B(_1167_),
    .Y(_0911_)
  );
  NOR _1773_ (
    .A(_0767_),
    .B(_1302_),
    .Y(_0912_)
  );
  NOR _1774_ (
    .A(_0912_),
    .B(_0911_),
    .Y(_0913_)
  );
  NAND _1775_ (
    .A(_0913_),
    .B(_0544_),
    .Y(_0914_)
  );
  NOR _1776_ (
    .A(_0914_),
    .B(_0910_),
    .Y(_0915_)
  );
  NOT _1777_ (
    .A(_0915_),
    .Y(_0916_)
  );
  NOR _1778_ (
    .A(_0916_),
    .B(_0909_),
    .Y(_0917_)
  );
  NOT _1779_ (
    .A(_0917_),
    .Y(_0918_)
  );
  NOR _1780_ (
    .A(_0918_),
    .B(_0903_),
    .Y(_0919_)
  );
  NAND _1781_ (
    .A(_0919_),
    .B(_0900_),
    .Y(_0920_)
  );
  NAND _1782_ (
    .A(_0920_),
    .B(_0895_),
    .Y(_0921_)
  );
  NOT _1783_ (
    .A(_0921_),
    .Y(_0685_)
  );
  NOR _1784_ (
    .A(_1232_),
    .B(_1209_),
    .Y(_0922_)
  );
  NAND _1785_ (
    .A(_0922_),
    .B(_0531_),
    .Y(_0923_)
  );
  NOR _1786_ (
    .A(_0922_),
    .B(_0531_),
    .Y(_0924_)
  );
  NOR _1787_ (
    .A(_0924_),
    .B(_0544_),
    .Y(_0925_)
  );
  NAND _1788_ (
    .A(_0925_),
    .B(_0923_),
    .Y(_0926_)
  );
  NOT _1789_ (
    .A(_0628_),
    .Y(_0927_)
  );
  NAND _1790_ (
    .A(_0564_),
    .B(_0562_),
    .Y(_0928_)
  );
  NOR _1791_ (
    .A(_0928_),
    .B(_0927_),
    .Y(_0929_)
  );
  NAND _1792_ (
    .A(_0928_),
    .B(_0927_),
    .Y(_0930_)
  );
  NAND _1793_ (
    .A(_0930_),
    .B(_0643_),
    .Y(_0931_)
  );
  NOR _1794_ (
    .A(_0931_),
    .B(_0929_),
    .Y(_0932_)
  );
  NOT _1795_ (
    .A(_0657_),
    .Y(_0933_)
  );
  NOT _1796_ (
    .A(_0659_),
    .Y(_0935_)
  );
  NOT _1797_ (
    .A(_0716_),
    .Y(_0936_)
  );
  NOR _1798_ (
    .A(_0936_),
    .B(_0713_),
    .Y(_0937_)
  );
  NOR _1799_ (
    .A(_0937_),
    .B(_0935_),
    .Y(_0938_)
  );
  NOT _1800_ (
    .A(_0938_),
    .Y(_0939_)
  );
  NAND _1801_ (
    .A(_0939_),
    .B(_0933_),
    .Y(_0940_)
  );
  NAND _1802_ (
    .A(_0940_),
    .B(_0662_),
    .Y(_0941_)
  );
  NOR _1803_ (
    .A(_0940_),
    .B(_0662_),
    .Y(_0942_)
  );
  NOR _1804_ (
    .A(_0942_),
    .B(_0733_),
    .Y(_0943_)
  );
  NAND _1805_ (
    .A(_0943_),
    .B(_0941_),
    .Y(_0944_)
  );
  NOT _1806_ (
    .A(_0748_),
    .Y(_0946_)
  );
  NOR _1807_ (
    .A(_0946_),
    .B(_1020_),
    .Y(_0947_)
  );
  NAND _1808_ (
    .A(_0750_),
    .B(_0757_),
    .Y(_0948_)
  );
  NOR _1809_ (
    .A(_0948_),
    .B(_0947_),
    .Y(_0949_)
  );
  NAND _1810_ (
    .A(_0769_),
    .B(_1242_),
    .Y(_0950_)
  );
  NOR _1811_ (
    .A(_0767_),
    .B(_1020_),
    .Y(_0951_)
  );
  NOR _1812_ (
    .A(_0848_),
    .B(_1221_),
    .Y(_0952_)
  );
  NOR _1813_ (
    .A(_0952_),
    .B(_0951_),
    .Y(_0953_)
  );
  NAND _1814_ (
    .A(_0953_),
    .B(_0950_),
    .Y(_0954_)
  );
  NOR _1815_ (
    .A(_0954_),
    .B(_0949_),
    .Y(_0955_)
  );
  NAND _1816_ (
    .A(_0955_),
    .B(_0944_),
    .Y(_0957_)
  );
  NOR _1817_ (
    .A(_0957_),
    .B(_0932_),
    .Y(_0958_)
  );
  NAND _1818_ (
    .A(_0958_),
    .B(_0926_),
    .Y(_0712_)
  );
  NOR _1819_ (
    .A(_0529_),
    .B(_1294_),
    .Y(_0959_)
  );
  NOR _1820_ (
    .A(_0959_),
    .B(_0813_),
    .Y(_0960_)
  );
  NOR _1821_ (
    .A(_0960_),
    .B(_0544_),
    .Y(_0961_)
  );
  NOT _1822_ (
    .A(_0961_),
    .Y(_0962_)
  );
  NOR _1823_ (
    .A(_0626_),
    .B(_0569_),
    .Y(_0963_)
  );
  NOT _1824_ (
    .A(_0963_),
    .Y(_0964_)
  );
  NAND _1825_ (
    .A(_0964_),
    .B(_0627_),
    .Y(_0965_)
  );
  NOR _1826_ (
    .A(_0965_),
    .B(_0830_),
    .Y(_0967_)
  );
  NOT _1827_ (
    .A(_0967_),
    .Y(_0968_)
  );
  NAND _1828_ (
    .A(_0937_),
    .B(_0935_),
    .Y(_0969_)
  );
  NAND _1829_ (
    .A(_0969_),
    .B(_0939_),
    .Y(_0970_)
  );
  NOR _1830_ (
    .A(_0970_),
    .B(_0733_),
    .Y(_0971_)
  );
  NOR _1831_ (
    .A(_0839_),
    .B(_1054_),
    .Y(_0972_)
  );
  NOR _1832_ (
    .A(_0946_),
    .B(_0878_),
    .Y(_0973_)
  );
  NOT _1833_ (
    .A(_0973_),
    .Y(_0974_)
  );
  NOR _1834_ (
    .A(_0974_),
    .B(_0972_),
    .Y(_0975_)
  );
  NOR _1835_ (
    .A(_0542_),
    .B(_1284_),
    .Y(_0976_)
  );
  NOR _1836_ (
    .A(_0976_),
    .B(_0543_),
    .Y(_0978_)
  );
  NOR _1837_ (
    .A(_0770_),
    .B(_1293_),
    .Y(_0979_)
  );
  NOR _1838_ (
    .A(_0767_),
    .B(_1054_),
    .Y(_0980_)
  );
  NOR _1839_ (
    .A(_0980_),
    .B(_0979_),
    .Y(_0981_)
  );
  NAND _1840_ (
    .A(_0981_),
    .B(_0978_),
    .Y(_0982_)
  );
  NOR _1841_ (
    .A(_0982_),
    .B(_0975_),
    .Y(_0983_)
  );
  NOT _1842_ (
    .A(_0983_),
    .Y(_0984_)
  );
  NOR _1843_ (
    .A(_0984_),
    .B(_0971_),
    .Y(_0985_)
  );
  NAND _1844_ (
    .A(_0985_),
    .B(_0968_),
    .Y(_0986_)
  );
  NAND _1845_ (
    .A(_0986_),
    .B(_0962_),
    .Y(_0987_)
  );
  NOT _1846_ (
    .A(_0987_),
    .Y(_0725_)
  );
  NOR _1847_ (
    .A(_0572_),
    .B(_0570_),
    .Y(_0989_)
  );
  NOR _1848_ (
    .A(_0989_),
    .B(_0624_),
    .Y(_0990_)
  );
  NAND _1849_ (
    .A(_0989_),
    .B(_0624_),
    .Y(_0991_)
  );
  NAND _1850_ (
    .A(_0991_),
    .B(_0643_),
    .Y(_0992_)
  );
  NOR _1851_ (
    .A(_0992_),
    .B(_0990_),
    .Y(_0993_)
  );
  NAND _1852_ (
    .A(_0711_),
    .B(_0837_),
    .Y(_0994_)
  );
  NAND _1853_ (
    .A(_0994_),
    .B(_0667_),
    .Y(_0995_)
  );
  NOR _1854_ (
    .A(_0994_),
    .B(_0667_),
    .Y(_0996_)
  );
  NOR _1855_ (
    .A(_0996_),
    .B(_0733_),
    .Y(_0997_)
  );
  NAND _1856_ (
    .A(_0997_),
    .B(_0995_),
    .Y(_0999_)
  );
  NOR _1857_ (
    .A(_0747_),
    .B(_1099_),
    .Y(_1000_)
  );
  NAND _1858_ (
    .A(_0840_),
    .B(_0757_),
    .Y(_1001_)
  );
  NOR _1859_ (
    .A(_1001_),
    .B(_1000_),
    .Y(_1002_)
  );
  NOT _1860_ (
    .A(_1301_),
    .Y(_1003_)
  );
  NOR _1861_ (
    .A(_0848_),
    .B(_1003_),
    .Y(_1004_)
  );
  NOR _1862_ (
    .A(_1004_),
    .B(_0543_),
    .Y(_1005_)
  );
  NOR _1863_ (
    .A(_0767_),
    .B(_1099_),
    .Y(_1006_)
  );
  NOR _1864_ (
    .A(_0770_),
    .B(_1296_),
    .Y(_1007_)
  );
  NOR _1865_ (
    .A(_1007_),
    .B(_1006_),
    .Y(_1008_)
  );
  NAND _1866_ (
    .A(_1008_),
    .B(_1005_),
    .Y(_1010_)
  );
  NOR _1867_ (
    .A(_1010_),
    .B(_1002_),
    .Y(_1011_)
  );
  NAND _1868_ (
    .A(_1011_),
    .B(_0999_),
    .Y(_1012_)
  );
  NOR _1869_ (
    .A(_1012_),
    .B(_0993_),
    .Y(_1013_)
  );
  NOR _1870_ (
    .A(_1296_),
    .B(_1301_),
    .Y(_1014_)
  );
  NOR _1871_ (
    .A(_1014_),
    .B(_0810_),
    .Y(_1015_)
  );
  NAND _1872_ (
    .A(_1014_),
    .B(_0810_),
    .Y(_1016_)
  );
  NAND _1873_ (
    .A(_1016_),
    .B(_0543_),
    .Y(_1017_)
  );
  NOR _1874_ (
    .A(_1017_),
    .B(_1015_),
    .Y(_1018_)
  );
  NOR _1875_ (
    .A(_1018_),
    .B(_1013_),
    .Y(_0745_)
  );
  NOR _1876_ (
    .A(_0525_),
    .B(_1308_),
    .Y(_1021_)
  );
  NOR _1877_ (
    .A(_1021_),
    .B(_0809_),
    .Y(_1022_)
  );
  NOR _1878_ (
    .A(_1022_),
    .B(_0544_),
    .Y(_1023_)
  );
  NOR _1879_ (
    .A(_0622_),
    .B(_0577_),
    .Y(_1024_)
  );
  NOT _1880_ (
    .A(_1024_),
    .Y(_1025_)
  );
  NAND _1881_ (
    .A(_1025_),
    .B(_0623_),
    .Y(_1026_)
  );
  NOR _1882_ (
    .A(_1026_),
    .B(_0830_),
    .Y(_1027_)
  );
  NOR _1883_ (
    .A(_0710_),
    .B(_0672_),
    .Y(_1028_)
  );
  NAND _1884_ (
    .A(_0734_),
    .B(_0711_),
    .Y(_1029_)
  );
  NOR _1885_ (
    .A(_1029_),
    .B(_1028_),
    .Y(_1030_)
  );
  NAND _1886_ (
    .A(_0838_),
    .B(_1304_),
    .Y(_1033_)
  );
  NOR _1887_ (
    .A(_0747_),
    .B(_0878_),
    .Y(_1034_)
  );
  NAND _1888_ (
    .A(_1034_),
    .B(_1033_),
    .Y(_1035_)
  );
  NOT _1889_ (
    .A(_1035_),
    .Y(_1036_)
  );
  NOR _1890_ (
    .A(_0542_),
    .B(_1306_),
    .Y(_1037_)
  );
  NOR _1891_ (
    .A(_1037_),
    .B(_0543_),
    .Y(_1038_)
  );
  NOR _1892_ (
    .A(_0770_),
    .B(_1307_),
    .Y(_1039_)
  );
  NOR _1893_ (
    .A(_0767_),
    .B(_1134_),
    .Y(_1040_)
  );
  NOR _1894_ (
    .A(_1040_),
    .B(_1039_),
    .Y(_1041_)
  );
  NAND _1895_ (
    .A(_1041_),
    .B(_1038_),
    .Y(_1042_)
  );
  NOR _1896_ (
    .A(_1042_),
    .B(_1036_),
    .Y(_1044_)
  );
  NOT _1897_ (
    .A(_1044_),
    .Y(_1045_)
  );
  NOR _1898_ (
    .A(_1045_),
    .B(_1030_),
    .Y(_1046_)
  );
  NOT _1899_ (
    .A(_1046_),
    .Y(_1047_)
  );
  NOR _1900_ (
    .A(_1047_),
    .B(_1027_),
    .Y(_1048_)
  );
  NOR _1901_ (
    .A(_1048_),
    .B(_1023_),
    .Y(_0765_)
  );
  NOT _1902_ (
    .A(_0620_),
    .Y(_1049_)
  );
  NAND _1903_ (
    .A(_0581_),
    .B(_0579_),
    .Y(_1050_)
  );
  NOR _1904_ (
    .A(_1050_),
    .B(_1049_),
    .Y(_1051_)
  );
  NAND _1905_ (
    .A(_1050_),
    .B(_1049_),
    .Y(_1052_)
  );
  NAND _1906_ (
    .A(_1052_),
    .B(_0643_),
    .Y(_1055_)
  );
  NOR _1907_ (
    .A(_1055_),
    .B(_1051_),
    .Y(_1056_)
  );
  NOT _1908_ (
    .A(_0708_),
    .Y(_1057_)
  );
  NAND _1909_ (
    .A(_1057_),
    .B(_0706_),
    .Y(_1058_)
  );
  NOR _1910_ (
    .A(_0704_),
    .B(_0673_),
    .Y(_1059_)
  );
  NAND _1911_ (
    .A(_1059_),
    .B(_1058_),
    .Y(_1060_)
  );
  NOR _1912_ (
    .A(_1059_),
    .B(_1058_),
    .Y(_1061_)
  );
  NOR _1913_ (
    .A(_1061_),
    .B(_0733_),
    .Y(_1062_)
  );
  NAND _1914_ (
    .A(_1062_),
    .B(_1060_),
    .Y(_1063_)
  );
  NOR _1915_ (
    .A(_0744_),
    .B(_0729_),
    .Y(_1064_)
  );
  NAND _1916_ (
    .A(_0838_),
    .B(_0757_),
    .Y(_1067_)
  );
  NOR _1917_ (
    .A(_1067_),
    .B(_1064_),
    .Y(_1068_)
  );
  NOT _1918_ (
    .A(_0463_),
    .Y(_1069_)
  );
  NOR _1919_ (
    .A(_0848_),
    .B(_1069_),
    .Y(_1070_)
  );
  NOR _1920_ (
    .A(_1070_),
    .B(_0543_),
    .Y(_1071_)
  );
  NOR _1921_ (
    .A(_0767_),
    .B(_0729_),
    .Y(_1072_)
  );
  NOR _1922_ (
    .A(_0770_),
    .B(_1309_),
    .Y(_1073_)
  );
  NOR _1923_ (
    .A(_1073_),
    .B(_1072_),
    .Y(_1074_)
  );
  NAND _1924_ (
    .A(_1074_),
    .B(_1071_),
    .Y(_1075_)
  );
  NOR _1925_ (
    .A(_1075_),
    .B(_1068_),
    .Y(_1076_)
  );
  NAND _1926_ (
    .A(_1076_),
    .B(_1063_),
    .Y(_1078_)
  );
  NOR _1927_ (
    .A(_1078_),
    .B(_1056_),
    .Y(_1079_)
  );
  NOR _1928_ (
    .A(_1309_),
    .B(_0463_),
    .Y(_1080_)
  );
  NOR _1929_ (
    .A(_1080_),
    .B(_0523_),
    .Y(_1081_)
  );
  NOT _1930_ (
    .A(_1080_),
    .Y(_1082_)
  );
  NOR _1931_ (
    .A(_1082_),
    .B(_0804_),
    .Y(_1083_)
  );
  NOR _1932_ (
    .A(_1083_),
    .B(_1081_),
    .Y(_1084_)
  );
  NOR _1933_ (
    .A(_1084_),
    .B(_0544_),
    .Y(_1085_)
  );
  NOR _1934_ (
    .A(_1085_),
    .B(_1079_),
    .Y(_0792_)
  );
  NOR _1935_ (
    .A(_0521_),
    .B(_0472_),
    .Y(_1086_)
  );
  NOR _1936_ (
    .A(_1086_),
    .B(_0803_),
    .Y(_1088_)
  );
  NOR _1937_ (
    .A(_1088_),
    .B(_0544_),
    .Y(_1089_)
  );
  NOR _1938_ (
    .A(_0618_),
    .B(_0585_),
    .Y(_1090_)
  );
  NOT _1939_ (
    .A(_1090_),
    .Y(_1091_)
  );
  NAND _1940_ (
    .A(_1091_),
    .B(_0619_),
    .Y(_1092_)
  );
  NOR _1941_ (
    .A(_1092_),
    .B(_0830_),
    .Y(_1093_)
  );
  NAND _1942_ (
    .A(_0703_),
    .B(_0677_),
    .Y(_1094_)
  );
  NOR _1943_ (
    .A(_0733_),
    .B(_0704_),
    .Y(_1095_)
  );
  NAND _1944_ (
    .A(_1095_),
    .B(_1094_),
    .Y(_1096_)
  );
  NOR _1945_ (
    .A(_0743_),
    .B(_0476_),
    .Y(_1097_)
  );
  NOR _1946_ (
    .A(_1097_),
    .B(_0762_),
    .Y(_1100_)
  );
  NOT _1947_ (
    .A(_0744_),
    .Y(_1101_)
  );
  NAND _1948_ (
    .A(_1101_),
    .B(_0757_),
    .Y(_1102_)
  );
  NOR _1949_ (
    .A(_1102_),
    .B(_1100_),
    .Y(_1103_)
  );
  NOR _1950_ (
    .A(_0770_),
    .B(_0470_),
    .Y(_1104_)
  );
  NOR _1951_ (
    .A(_1104_),
    .B(_0543_),
    .Y(_1105_)
  );
  NOR _1952_ (
    .A(_0767_),
    .B(_0762_),
    .Y(_1106_)
  );
  NOR _1953_ (
    .A(_0848_),
    .B(_0468_),
    .Y(_1107_)
  );
  NOR _1954_ (
    .A(_1107_),
    .B(_1106_),
    .Y(_1108_)
  );
  NAND _1955_ (
    .A(_1108_),
    .B(_1105_),
    .Y(_1109_)
  );
  NOR _1956_ (
    .A(_1109_),
    .B(_1103_),
    .Y(_1113_)
  );
  NAND _1957_ (
    .A(_1113_),
    .B(_1096_),
    .Y(_1114_)
  );
  NOR _1958_ (
    .A(_1114_),
    .B(_1093_),
    .Y(_1115_)
  );
  NOR _1959_ (
    .A(_1115_),
    .B(_1089_),
    .Y(_0805_)
  );
  NOR _1960_ (
    .A(_0473_),
    .B(_0477_),
    .Y(_1116_)
  );
  NOT _1961_ (
    .A(_1116_),
    .Y(_1117_)
  );
  NAND _1962_ (
    .A(_1117_),
    .B(_0519_),
    .Y(_1118_)
  );
  NAND _1963_ (
    .A(_1116_),
    .B(_0800_),
    .Y(_1119_)
  );
  NAND _1964_ (
    .A(_1119_),
    .B(_1118_),
    .Y(_1120_)
  );
  NAND _1965_ (
    .A(_1120_),
    .B(_0543_),
    .Y(_1121_)
  );
  NOR _1966_ (
    .A(_0588_),
    .B(_0586_),
    .Y(_1123_)
  );
  NAND _1967_ (
    .A(_1123_),
    .B(_0616_),
    .Y(_1124_)
  );
  NOT _1968_ (
    .A(_0616_),
    .Y(_1125_)
  );
  NOT _1969_ (
    .A(_1123_),
    .Y(_1126_)
  );
  NAND _1970_ (
    .A(_1126_),
    .B(_1125_),
    .Y(_1127_)
  );
  NAND _1971_ (
    .A(_1127_),
    .B(_1124_),
    .Y(_1128_)
  );
  NOR _1972_ (
    .A(_1128_),
    .B(_0830_),
    .Y(_1129_)
  );
  NOT _1973_ (
    .A(_0679_),
    .Y(_1130_)
  );
  NAND _1974_ (
    .A(_1130_),
    .B(_0736_),
    .Y(_1131_)
  );
  NAND _1975_ (
    .A(_1131_),
    .B(_0701_),
    .Y(_1132_)
  );
  NOR _1976_ (
    .A(_1131_),
    .B(_0701_),
    .Y(_1135_)
  );
  NOR _1977_ (
    .A(_1135_),
    .B(_0733_),
    .Y(_1136_)
  );
  NAND _1978_ (
    .A(_1136_),
    .B(_1132_),
    .Y(_1137_)
  );
  NAND _1979_ (
    .A(_0743_),
    .B(_0476_),
    .Y(_1138_)
  );
  NAND _1980_ (
    .A(_1138_),
    .B(_0757_),
    .Y(_1139_)
  );
  NOR _1981_ (
    .A(_1139_),
    .B(_1097_),
    .Y(_1140_)
  );
  NAND _1982_ (
    .A(_0763_),
    .B(_0477_),
    .Y(_1141_)
  );
  NOR _1983_ (
    .A(_0770_),
    .B(_0473_),
    .Y(_1142_)
  );
  NOR _1984_ (
    .A(_0767_),
    .B(_0807_),
    .Y(_1143_)
  );
  NOR _1985_ (
    .A(_1143_),
    .B(_1142_),
    .Y(_1144_)
  );
  NAND _1986_ (
    .A(_1144_),
    .B(_1141_),
    .Y(_1147_)
  );
  NOR _1987_ (
    .A(_1147_),
    .B(_1140_),
    .Y(_1148_)
  );
  NAND _1988_ (
    .A(_1148_),
    .B(_1137_),
    .Y(_1149_)
  );
  NOR _1989_ (
    .A(_1149_),
    .B(_1129_),
    .Y(_1150_)
  );
  NAND _1990_ (
    .A(_1150_),
    .B(_1121_),
    .Y(_0822_)
  );
  NOR _1991_ (
    .A(_0517_),
    .B(_0483_),
    .Y(_1151_)
  );
  NOR _1992_ (
    .A(_1151_),
    .B(_0799_),
    .Y(_1152_)
  );
  NOR _1993_ (
    .A(_1152_),
    .B(_0544_),
    .Y(_1153_)
  );
  NOR _1994_ (
    .A(_0614_),
    .B(_0594_),
    .Y(_1154_)
  );
  NOT _1995_ (
    .A(_0615_),
    .Y(_1155_)
  );
  NOR _1996_ (
    .A(_0830_),
    .B(_1155_),
    .Y(_1157_)
  );
  NOT _1997_ (
    .A(_1157_),
    .Y(_1158_)
  );
  NOR _1998_ (
    .A(_1158_),
    .B(_1154_),
    .Y(_1159_)
  );
  NAND _1999_ (
    .A(_0699_),
    .B(_0683_),
    .Y(_1160_)
  );
  NOR _2000_ (
    .A(_0733_),
    .B(_0700_),
    .Y(_1161_)
  );
  NAND _2001_ (
    .A(_1161_),
    .B(_1160_),
    .Y(_1162_)
  );
  NOR _2002_ (
    .A(_0741_),
    .B(_0486_),
    .Y(_1163_)
  );
  NOR _2003_ (
    .A(_1163_),
    .B(_0841_),
    .Y(_1164_)
  );
  NAND _2004_ (
    .A(_0743_),
    .B(_0757_),
    .Y(_1165_)
  );
  NOR _2005_ (
    .A(_1165_),
    .B(_1164_),
    .Y(_1166_)
  );
  NOR _2006_ (
    .A(_0542_),
    .B(_0481_),
    .Y(_1168_)
  );
  NOR _2007_ (
    .A(_1168_),
    .B(_0543_),
    .Y(_1169_)
  );
  NOR _2008_ (
    .A(_0770_),
    .B(_0482_),
    .Y(_1170_)
  );
  NOR _2009_ (
    .A(_0767_),
    .B(_0841_),
    .Y(_1171_)
  );
  NOR _2010_ (
    .A(_1171_),
    .B(_1170_),
    .Y(_1172_)
  );
  NAND _2011_ (
    .A(_1172_),
    .B(_1169_),
    .Y(_1173_)
  );
  NOR _2012_ (
    .A(_1173_),
    .B(_1166_),
    .Y(_1174_)
  );
  NAND _2013_ (
    .A(_1174_),
    .B(_1162_),
    .Y(_1175_)
  );
  NOR _2014_ (
    .A(_1175_),
    .B(_1159_),
    .Y(_1176_)
  );
  NOR _2015_ (
    .A(_1176_),
    .B(_1153_),
    .Y(_0836_)
  );
  NOR _2016_ (
    .A(_0489_),
    .B(_0487_),
    .Y(_1178_)
  );
  NAND _2017_ (
    .A(_1178_),
    .B(_0796_),
    .Y(_1179_)
  );
  NOT _2018_ (
    .A(_1178_),
    .Y(_1180_)
  );
  NAND _2019_ (
    .A(_1180_),
    .B(_0514_),
    .Y(_1181_)
  );
  NAND _2020_ (
    .A(_1181_),
    .B(_1179_),
    .Y(_1182_)
  );
  NAND _2021_ (
    .A(_1182_),
    .B(_0543_),
    .Y(_1183_)
  );
  NOR _2022_ (
    .A(_0612_),
    .B(_0610_),
    .Y(_1184_)
  );
  NAND _2023_ (
    .A(_0643_),
    .B(_0613_),
    .Y(_1185_)
  );
  NOR _2024_ (
    .A(_1185_),
    .B(_1184_),
    .Y(_1186_)
  );
  NOR _2025_ (
    .A(_0686_),
    .B(_0684_),
    .Y(_1187_)
  );
  NAND _2026_ (
    .A(_1187_),
    .B(_0696_),
    .Y(_1189_)
  );
  NOR _2027_ (
    .A(_1187_),
    .B(_0696_),
    .Y(_1190_)
  );
  NOR _2028_ (
    .A(_1190_),
    .B(_0733_),
    .Y(_1191_)
  );
  NAND _2029_ (
    .A(_1191_),
    .B(_1189_),
    .Y(_1192_)
  );
  NAND _2030_ (
    .A(_0741_),
    .B(_0486_),
    .Y(_1193_)
  );
  NAND _2031_ (
    .A(_1193_),
    .B(_0757_),
    .Y(_1194_)
  );
  NOR _2032_ (
    .A(_1194_),
    .B(_1163_),
    .Y(_1195_)
  );
  NAND _2033_ (
    .A(_0769_),
    .B(_0490_),
    .Y(_1196_)
  );
  NOR _2034_ (
    .A(_0767_),
    .B(_0568_),
    .Y(_1197_)
  );
  NOR _2035_ (
    .A(_0848_),
    .B(_0488_),
    .Y(_1198_)
  );
  NOR _2036_ (
    .A(_1198_),
    .B(_1197_),
    .Y(_1200_)
  );
  NAND _2037_ (
    .A(_1200_),
    .B(_1196_),
    .Y(_1201_)
  );
  NOR _2038_ (
    .A(_1201_),
    .B(_1195_),
    .Y(_1202_)
  );
  NAND _2039_ (
    .A(_1202_),
    .B(_1192_),
    .Y(_1203_)
  );
  NOR _2040_ (
    .A(_1203_),
    .B(_1186_),
    .Y(_1204_)
  );
  NAND _2041_ (
    .A(_1204_),
    .B(_1183_),
    .Y(_0856_)
  );
  NOR _2042_ (
    .A(_0512_),
    .B(_0496_),
    .Y(_1205_)
  );
  NOR _2043_ (
    .A(_1205_),
    .B(_0794_),
    .Y(_1206_)
  );
  NOR _2044_ (
    .A(_1206_),
    .B(_0544_),
    .Y(_1207_)
  );
  NOR _2045_ (
    .A(_0608_),
    .B(_0606_),
    .Y(_1208_)
  );
  NOT _2046_ (
    .A(_1208_),
    .Y(_1210_)
  );
  NAND _2047_ (
    .A(_1210_),
    .B(_0609_),
    .Y(_1211_)
  );
  NOR _2048_ (
    .A(_1211_),
    .B(_0830_),
    .Y(_1212_)
  );
  NAND _2049_ (
    .A(_0693_),
    .B(_0690_),
    .Y(_1213_)
  );
  NAND _2050_ (
    .A(_1213_),
    .B(_0734_),
    .Y(_1214_)
  );
  NOR _2051_ (
    .A(_1214_),
    .B(_0694_),
    .Y(_1215_)
  );
  NOR _2052_ (
    .A(_0738_),
    .B(_0600_),
    .Y(_1216_)
  );
  NOT _2053_ (
    .A(_1216_),
    .Y(_1217_)
  );
  NAND _2054_ (
    .A(_1217_),
    .B(_0741_),
    .Y(_1218_)
  );
  NOR _2055_ (
    .A(_1218_),
    .B(_0878_),
    .Y(_1219_)
  );
  NOR _2056_ (
    .A(_0767_),
    .B(_0600_),
    .Y(_1222_)
  );
  NOR _2057_ (
    .A(_1222_),
    .B(_0543_),
    .Y(_1223_)
  );
  NOR _2058_ (
    .A(_0770_),
    .B(_0495_),
    .Y(_1224_)
  );
  NOR _2059_ (
    .A(_0848_),
    .B(_0494_),
    .Y(_1225_)
  );
  NOR _2060_ (
    .A(_1225_),
    .B(_1224_),
    .Y(_1226_)
  );
  NAND _2061_ (
    .A(_1226_),
    .B(_1223_),
    .Y(_1227_)
  );
  NOR _2062_ (
    .A(_1227_),
    .B(_1219_),
    .Y(_1228_)
  );
  NOT _2063_ (
    .A(_1228_),
    .Y(_1229_)
  );
  NOR _2064_ (
    .A(_1229_),
    .B(_1215_),
    .Y(_1230_)
  );
  NOT _2065_ (
    .A(_1230_),
    .Y(_1231_)
  );
  NOR _2066_ (
    .A(_1231_),
    .B(_1212_),
    .Y(_1233_)
  );
  NOR _2067_ (
    .A(_1233_),
    .B(_1207_),
    .Y(_0867_)
  );
  NOR _2068_ (
    .A(_0510_),
    .B(_0508_),
    .Y(_1234_)
  );
  NOR _2069_ (
    .A(_1234_),
    .B(_0791_),
    .Y(_1235_)
  );
  NOR _2070_ (
    .A(_1235_),
    .B(_0544_),
    .Y(_1236_)
  );
  NOR _2071_ (
    .A(_0600_),
    .B(_1220_),
    .Y(_1237_)
  );
  NOR _2072_ (
    .A(_1237_),
    .B(_0692_),
    .Y(_1238_)
  );
  NOR _2073_ (
    .A(_1238_),
    .B(_0740_),
    .Y(_1239_)
  );
  NOR _2074_ (
    .A(_1239_),
    .B(_0733_),
    .Y(_1240_)
  );
  NOR _2075_ (
    .A(_0767_),
    .B(_1220_),
    .Y(_1241_)
  );
  NOR _2076_ (
    .A(_0770_),
    .B(_0509_),
    .Y(_1243_)
  );
  NOR _2077_ (
    .A(_1243_),
    .B(_1241_),
    .Y(_1244_)
  );
  NOR _2078_ (
    .A(_0604_),
    .B(_0602_),
    .Y(_1245_)
  );
  NAND _2079_ (
    .A(_0643_),
    .B(_0605_),
    .Y(_1246_)
  );
  NOR _2080_ (
    .A(_1246_),
    .B(_1245_),
    .Y(_1247_)
  );
  NAND _2081_ (
    .A(_0503_),
    .B(_0498_),
    .Y(_1248_)
  );
  NAND _2082_ (
    .A(_1248_),
    .B(_0739_),
    .Y(_1249_)
  );
  NOR _2083_ (
    .A(_1249_),
    .B(_0878_),
    .Y(_1250_)
  );
  NOR _2084_ (
    .A(_1250_),
    .B(_0543_),
    .Y(_1251_)
  );
  NAND _2085_ (
    .A(_0763_),
    .B(_0499_),
    .Y(_1252_)
  );
  NAND _2086_ (
    .A(_1252_),
    .B(_1251_),
    .Y(_1254_)
  );
  NOR _2087_ (
    .A(_1254_),
    .B(_1247_),
    .Y(_1255_)
  );
  NAND _2088_ (
    .A(_1255_),
    .B(_1244_),
    .Y(_1256_)
  );
  NOR _2089_ (
    .A(_1256_),
    .B(_1240_),
    .Y(_1257_)
  );
  NOR _2090_ (
    .A(_1257_),
    .B(_1236_),
    .Y(_0880_)
  );
  NOR _2091_ (
    .A(_0485_),
    .B(_1111_),
    .Y(_1258_)
  );
  NOR _2092_ (
    .A(_1258_),
    .B(_0602_),
    .Y(_1259_)
  );
  NAND _2093_ (
    .A(_1259_),
    .B(_0643_),
    .Y(_1260_)
  );
  NOR _2094_ (
    .A(_0848_),
    .B(_0501_),
    .Y(_1261_)
  );
  NOR _2095_ (
    .A(_1249_),
    .B(_0733_),
    .Y(_1262_)
  );
  NOR _2096_ (
    .A(_1262_),
    .B(_1261_),
    .Y(_1264_)
  );
  NAND _2097_ (
    .A(_1264_),
    .B(_1260_),
    .Y(_1265_)
  );
  NAND _2098_ (
    .A(_0755_),
    .B(_0503_),
    .Y(_1266_)
  );
  NAND _2099_ (
    .A(_0769_),
    .B(_0786_),
    .Y(_1267_)
  );
  NAND _2100_ (
    .A(_1267_),
    .B(_1266_),
    .Y(_1268_)
  );
  NOR _2101_ (
    .A(_1268_),
    .B(_1265_),
    .Y(_1269_)
  );
  NOR _2102_ (
    .A(_0506_),
    .B(_0516_),
    .Y(_1270_)
  );
  NOR _2103_ (
    .A(_1270_),
    .B(_0788_),
    .Y(_1271_)
  );
  NAND _2104_ (
    .A(_1271_),
    .B(_0543_),
    .Y(_1272_)
  );
  NAND _2105_ (
    .A(_1272_),
    .B(_1269_),
    .Y(_0890_)
  );
  NOT _2106_ (
    .A(_0765_),
    .Y(_1274_)
  );
  NOT _2107_ (
    .A(_0805_),
    .Y(_1275_)
  );
  NOT _2108_ (
    .A(_0836_),
    .Y(_1276_)
  );
  NOT _2109_ (
    .A(_0867_),
    .Y(_1277_)
  );
  NOR _2110_ (
    .A(_0890_),
    .B(_0880_),
    .Y(_1278_)
  );
  NAND _2111_ (
    .A(_1278_),
    .B(_1277_),
    .Y(_1279_)
  );
  NOR _2112_ (
    .A(_1279_),
    .B(_0856_),
    .Y(_1280_)
  );
  NAND _2113_ (
    .A(_1280_),
    .B(_1276_),
    .Y(_1281_)
  );
  NOR _2114_ (
    .A(_1281_),
    .B(_0822_),
    .Y(_1282_)
  );
  NAND _2115_ (
    .A(_1282_),
    .B(_1275_),
    .Y(_1283_)
  );
  NOR _2116_ (
    .A(_1283_),
    .B(_0792_),
    .Y(_1285_)
  );
  NAND _2117_ (
    .A(_1285_),
    .B(_1274_),
    .Y(_1286_)
  );
  NOR _2118_ (
    .A(_1286_),
    .B(_0745_),
    .Y(_1287_)
  );
  NAND _2119_ (
    .A(_1287_),
    .B(_0987_),
    .Y(_1288_)
  );
  NOR _2120_ (
    .A(_1288_),
    .B(_0712_),
    .Y(_1289_)
  );
  NAND _2121_ (
    .A(_1289_),
    .B(_0921_),
    .Y(_1290_)
  );
  NOR _2122_ (
    .A(_1290_),
    .B(_0669_),
    .Y(_1291_)
  );
  NAND _2123_ (
    .A(_1291_),
    .B(_0860_),
    .Y(_1292_)
  );
  NOR _2124_ (
    .A(_1292_),
    .B(_0638_),
    .Y(_0905_)
  );
  assign outF[15] = neg;
  assign _0459_ = inN[15];
  assign _0460_ = inM[15];
  assign _0674_ = inN[14];
  assign _0783_ = inM[14];
  assign _1111_ = inN[1];
  assign _1220_ = inM[1];
  assign _0474_ = inN[0];
  assign _0485_ = inM[0];
  assign _0516_ = inC;
  assign _0557_ = inN[3];
  assign _0568_ = inM[3];
  assign _0589_ = inN[2];
  assign _0600_ = inM[2];
  assign _0717_ = inN[7];
  assign _0729_ = inM[7];
  assign _0751_ = inN[6];
  assign _0762_ = inM[6];
  assign _0795_ = inN[5];
  assign _0807_ = inM[5];
  assign _0829_ = inN[4];
  assign _0841_ = inM[4];
  assign _1009_ = inN[11];
  assign _1020_ = inM[11];
  assign _1043_ = inN[10];
  assign _1054_ = inM[10];
  assign _1087_ = inN[9];
  assign _1099_ = inM[9];
  assign _1122_ = inN[8];
  assign _1134_ = inM[8];
  assign _1295_ = inN[13];
  assign _1297_ = inM[13];
  assign _1300_ = inN[12];
  assign _1302_ = inM[12];
  assign _0466_ = opc[2];
  assign _0469_ = opc[1];
  assign _0471_ = opc[0];
  assign neg = _0638_;
  assign outF[14] = _0650_;
  assign outF[13] = _0669_;
  assign outF[12] = _0685_;
  assign outF[11] = _0712_;
  assign outF[10] = _0725_;
  assign outF[9] = _0745_;
  assign outF[8] = _0765_;
  assign outF[7] = _0792_;
  assign outF[6] = _0805_;
  assign outF[5] = _0822_;
  assign outF[4] = _0836_;
  assign outF[3] = _0856_;
  assign outF[2] = _0867_;
  assign outF[1] = _0880_;
  assign outF[0] = _0890_;
  assign zer = _0905_;
endmodule
