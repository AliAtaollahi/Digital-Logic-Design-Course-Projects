`timescale 1ns/1ns
module mux2_to_1 (input a,b,s,en,output w);
	wire i,j;
	notif1 #(14,18,16) n1(i,a,j);
	notif1 #(14,18,16) n2(i,b,s);
	not #(7,9) n3(j,s);
	notif1 #(14,18,16) n4(w,i,en);
endmodule
module D_latch(input d,clk,en,output q);
	mux2_to_1 mx(q,d,clk,en,q);
endmodule
module register8withDlatch(input serIn,clk,en,output [7:0] po);
	wire [8:0] d;
	assign d[8]=serIn;
	genvar k;
	generate
		for(k=8;k>0;k=k-1) begin : registerGates
			D_latch dd(d[k],clk,en,d[k-1]);
		end
	endgenerate
	assign po=d[7:0];
endmodule