`timescale 1ns/1ns
module mult (input [15:0] a,b,output [31:0] w);
	assign w=a*b;
endmodule
